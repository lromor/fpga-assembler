module top (
    output wire ja0,
    input  wire ja1
);
  assign ja0 = ja1;
endmodule
